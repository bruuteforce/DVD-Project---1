*cfr3-BandAn -- Indipendent signal generators and Vdd power supply
*(AandB)n for all combinations of input.

.INCLUDE 45nm_HP.pm
.OPTIONS GMIN=1e-020 ABSTOL=1e-018

*Definition 
.PARAM Lmin=45n
.PARAM Ldiff=90n
.PARAM Wmin=45n

Vdd 	vgen 	0 
Va 	A 	0 	
Vb 	B 	0 
Vbody1 b1	0	1.1
Vbody2	b2	0	1.1

Mn1 	SD1 	A 	0 		b2 	pmos W={Wmin} L={Lmin}
Mn2 	vgen 	B 	SD1 	b1 	pmos W={Wmin} L={Lmin} 

.TEMP 25
.CONTROL
echo "AandBn Stack" > AandBp.txt
let Ldiff=90n
foreach Vddbasic 1.1
  echo Vdd basic = $Vddbasic
   alter Vdd = $Vddbasic
	foreach width 45n
	echo Wmin=$width
			foreach input 0 $Vddbasic
		 	alter Va = $input
 	        			foreach input 0 $Vddbasic
					 alter Vb = $input
			        *if not(@Vdd[DC] & @Va[DC] & @Vb[DC] )
	 	echo DC Analysis at 25C          			
		dc TEMP 25 90 70
		print V(SD1) V(vgen) V(A) V(B) >> AandBp.txt
			   
			        end
			    end	
	    end
	end	
   
.ENDC
.END
