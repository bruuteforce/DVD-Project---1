*cfr3-BandAn -- Indipendent signal generators and Vdd power supply
*(AandB)n for all combinations of input.

.INCLUDE ../model/45nm_HP.pm
.OPTIONS GMIN=1e-020 ABSTOL=1e-018

*Definition 
.PARAM Lmin=45n
.PARAM Ldiff=90n
.PARAM Wmin=45n

Vdd 	vgen 	0 
Va 	A 	0 	
Vb 	B 	0 

Mn1 	SD1 	A 	0 		0 	nmos W={Wmin} L={Lmin}
Mn2 	vgen 	B 	SD1 	0 	nmos W={Wmin} L={Lmin} 

.TEMP 25

.CONTROL
echo "AandBn Stack" > AandBn.txt
let Ldiff=90n
foreach Vddbasic 1.1
  echo Vdd basic = $Vddbasic
   alter Vdd = $Vddbasic
	foreach width 45n

	echo
	echo
	echo Wmin=$width

			foreach input 0 $Vddbasic
		 	alter Va = $input
 	        			foreach input 0 $Vddbasic
					 alter Vb = $input
			        *if not(@Vdd[DC] & @Va[DC] & @Vb[DC] )
		

	 	echo DC Analysis at 25C
		            			
		dc TEMP 25 90 70
		print V(SD1) ((V(A)*(I(Va))+V(B)*(I(Vb))+V(vgen)*(I(Vdd)))) V(vgen) V(A) V(B) >> AandBn.txt
			   
			        end
			    end	
	    end
	end	
   
.ENDC
.END
