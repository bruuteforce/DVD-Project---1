*NMOS ON Condition

.INCLUDE 45nm_HP.pm

.PARAM Lmin=45n
.PARAM Wmin=45n
.PARAM Ldiff=90n
	
Mn drain gate source body nmos W={Wmin} L={Lmin} AS={Wmin*Ldiff} AD={Wmin*Ldiff} PS={2*(Ldiff+Wmin)} PD={2*(Ldiff+Wmin)}
Vd 	drain	d1		0
Vg 	gate	g1		0
Vs 	source	s1	  0
Vb 	body	0		0
Vdd 	d1	0		0
Vgg  g1  0  1.1
Vss  s1  0  0
.TEMP 25
.CONTROL
echo "NMOS ON Condition" > NMOS_on.txt
let voltage = 0
while voltage le 1.1125
  let voltage1 = 0
  alter Vss = 0
  while voltage1 le 1.1125
    dc TEMP 25 50 30
    print V(drain) V(gate) V(source) V(body) I(Vd) I(Vg) I(Vs) I(Vb) >> NMOS_on.txt
    let voltage1 = voltage1 + 0.025
    alter Vss = voltage1
  end
  let voltage = voltage + 0.025
  alter Vdd = voltage
end
.ENDC
.END